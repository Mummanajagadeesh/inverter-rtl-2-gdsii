// This is the unpowered netlist.
module inverter (in,
    out);
 input in;
 output out;

 wire net1;
 wire net2;

 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__inv_2 _0_ (.A(net1),
    .Y(net2));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 output2 (.A(net2),
    .X(out));
endmodule

