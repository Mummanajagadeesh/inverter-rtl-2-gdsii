VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO inverter
  CLASS BLOCK ;
  FOREIGN inverter ;
  ORIGIN 0.000 0.000 ;
  SIZE 34.500 BY 57.120 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 46.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 46.480 ;
    END
  END VPWR
  PIN in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 53.120 32.570 57.120 ;
    END
  END in
  PIN out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END out
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 28.980 46.325 ;
      LAYER met1 ;
        RECT 0.070 10.640 32.590 46.480 ;
      LAYER met2 ;
        RECT 0.100 52.840 32.010 53.120 ;
        RECT 0.100 4.280 32.560 52.840 ;
        RECT 0.650 4.000 32.560 4.280 ;
      LAYER met3 ;
        RECT 9.730 10.715 14.610 46.405 ;
  END
END inverter
END LIBRARY

