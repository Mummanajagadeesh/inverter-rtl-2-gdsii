magic
tech sky130A
magscale 1 2
timestamp 1758435569
<< checkpaint >>
rect -1298 -1860 2034 2452
rect 5220 -548 8920 652
rect 5220 -1748 10062 -548
rect 5220 -2948 10652 -1748
rect 5220 -3660 11426 -2948
rect 6362 -4148 11426 -3660
rect 6362 -4860 12568 -4148
rect 7504 -5348 12568 -4860
rect 7504 -6060 13710 -5348
rect 8094 -6548 13710 -6060
rect 8094 -7260 14300 -6548
rect 8868 -7748 14300 -7260
rect 8868 -8460 15442 -7748
rect 10010 -8948 15442 -8460
rect 10010 -9660 15642 -8948
rect 11152 -10148 15642 -9660
rect 11152 -10860 15956 -10148
rect 11742 -11348 15956 -10860
rect 11742 -12060 17098 -11348
rect 12884 -12548 17098 -12060
rect 12884 -13260 17412 -12548
rect 13084 -13748 17412 -13260
rect 13084 -14460 17612 -13748
rect 13398 -14948 17612 -14460
rect 13398 -15660 17926 -14948
rect 14540 -16148 17926 -15660
rect 14540 -16860 19068 -16148
rect 14854 -17348 19068 -16860
rect 14854 -18060 19382 -17348
rect 15054 -18548 19382 -18060
rect 15054 -19260 19582 -18548
rect 15368 -19748 19582 -19260
rect 15368 -20460 19896 -19748
rect 16510 -20948 19896 -20460
rect 16510 -21660 20096 -20948
rect 16824 -22148 20096 -21660
rect 16824 -22860 21238 -22148
rect 17024 -23348 21238 -22860
rect 17024 -24060 22380 -23348
rect 17338 -24548 22380 -24060
rect 17338 -25260 23154 -24548
rect 17538 -25748 23154 -25260
rect 17538 -26460 23468 -25748
rect 18680 -26948 23468 -26460
rect 18680 -27660 23668 -26948
rect 19822 -28148 23668 -27660
rect 19822 -28860 24810 -28148
rect 20596 -29348 24810 -28860
rect 20596 -30060 25400 -29348
rect 20910 -30548 25400 -30060
rect 20910 -31260 26542 -30548
rect 21110 -31748 26542 -31260
rect 21110 -32460 26856 -31748
rect 22252 -32948 26856 -32460
rect 22252 -33660 27998 -32948
rect 22842 -34148 27998 -33660
rect 22842 -34860 28198 -34148
rect 23984 -35348 28198 -34860
rect 23984 -36060 28512 -35348
rect 24298 -36548 28512 -36060
rect 24298 -37260 29654 -36548
rect 25440 -37748 29654 -37260
rect 25440 -38460 30796 -37748
rect 25640 -38948 30796 -38460
rect 25640 -39660 31110 -38948
rect 25954 -40860 31110 -39660
rect 27096 -40948 31110 -40860
rect 27096 -42060 31424 -40948
rect 28238 -42148 31424 -42060
rect 28238 -43348 32198 -42148
rect 28238 -44060 33340 -43348
rect 28552 -44548 33340 -44060
rect 28552 -45260 33654 -44548
rect 28866 -45748 33654 -45260
rect 28866 -46460 34244 -45748
rect 29640 -46948 34244 -46460
rect 29640 -47660 34558 -46948
rect 30782 -48148 34558 -47660
rect 30782 -48860 35700 -48148
rect 31096 -49348 35700 -48860
rect 31096 -50060 36842 -49348
rect 31686 -50548 36842 -50060
rect 31686 -51260 37432 -50548
rect 32000 -51748 37432 -51260
rect 32000 -52460 37632 -51748
rect 33142 -52948 37632 -52460
rect 33142 -53348 37832 -52948
rect 33142 -53660 38974 -53348
rect 34284 -54548 38974 -53660
rect 34284 -54860 40116 -54548
rect 34874 -55748 40116 -54860
rect 34874 -56060 40316 -55748
rect 35074 -56148 40316 -56060
rect 35074 -56460 40516 -56148
rect 35274 -56548 40516 -56460
rect 35274 -57660 41658 -56548
rect 36416 -57748 41658 -57660
rect 36416 -58860 41858 -57748
rect 37558 -58948 41858 -58860
rect 37558 -59260 42058 -58948
rect 37758 -59660 42058 -59260
rect 37958 -60148 42058 -59660
rect 37958 -60860 42832 -60148
rect 39100 -61348 42832 -60860
rect 39100 -62060 43146 -61348
rect 39300 -63260 43146 -62060
rect 39500 -63348 43146 -63260
rect 39500 -64460 44288 -63348
rect 40274 -64548 44288 -64460
rect 40274 -65748 44488 -64548
rect 40274 -66460 45630 -65748
rect 40588 -66948 45630 -66460
rect 40588 -67660 46772 -66948
rect 41730 -68148 46772 -67660
rect 41730 -68860 46972 -68148
rect 41930 -69348 46972 -68860
rect 41930 -70060 48114 -69348
rect 43072 -70548 48114 -70060
rect 43072 -71260 49256 -70548
rect 44214 -71748 49256 -71260
rect 44214 -72460 49456 -71748
rect 44414 -72948 49456 -72460
rect 44414 -73660 50230 -72948
rect 45556 -74148 50230 -73660
rect 45556 -74860 50636 -74148
rect 46698 -75348 50636 -74860
rect 46698 -76060 51778 -75348
rect 46898 -76548 51778 -76060
rect 46898 -77260 52092 -76548
rect 47672 -77748 52092 -77260
rect 47672 -78148 52292 -77748
rect 47672 -78460 52606 -78148
rect 48078 -79348 52606 -78460
rect 48078 -79660 53748 -79348
rect 49220 -80548 53748 -79660
rect 49220 -80860 54062 -80548
rect 49534 -81260 54062 -80860
rect 49734 -81748 54062 -81260
rect 49734 -82460 55204 -81748
rect 50048 -82948 55204 -82460
rect 50048 -83660 55794 -82948
rect 51190 -84148 55794 -83660
rect 51190 -84548 55994 -84148
rect 51190 -84860 56308 -84548
rect 51504 -85748 56308 -84860
rect 51504 -86060 56622 -85748
rect 52646 -86948 56622 -86060
rect 52646 -87260 56822 -86948
rect 53236 -87348 56822 -87260
rect 53236 -87660 57136 -87348
rect 53436 -88548 57136 -87660
rect 53436 -88860 57726 -88548
rect 53750 -89748 57726 -88860
rect 53750 -90060 58040 -89748
rect 54064 -90460 58040 -90060
rect 54264 -90948 58040 -90460
rect 54264 -91660 58630 -90948
rect 54578 -92148 58630 -91660
rect 54578 -92860 58944 -92148
rect 55168 -93348 58944 -92860
rect 55168 -94060 60086 -93348
rect 55482 -94548 60086 -94060
rect 55482 -94948 60286 -94548
rect 55482 -95260 60600 -94948
rect 56072 -96148 60600 -95260
rect 56072 -96460 60914 -96148
rect 56386 -97348 60914 -96460
rect 56386 -97660 61228 -97348
rect 57528 -98060 61228 -97660
rect 57728 -98548 61228 -98060
rect 57728 -99260 61542 -98548
rect 58042 -99748 61542 -99260
rect 58042 -100460 62684 -99748
rect 58356 -100948 62684 -100460
rect 58356 -101660 63274 -100948
rect 58670 -102860 63274 -101660
rect 58984 -102948 63274 -102860
rect 58984 -104060 64416 -102948
rect 60126 -104148 64416 -104060
rect 60126 -105348 64730 -104148
rect 60126 -106060 64930 -105348
rect 60716 -106548 64930 -106060
rect 60716 -107260 65244 -106548
rect 61858 -107748 65244 -107260
rect 61858 -108460 65444 -107748
rect 62172 -108948 65444 -108460
rect 62172 -109660 65644 -108948
rect 62372 -110148 65644 -109660
rect 62372 -110860 65844 -110148
rect 62686 -111348 65844 -110860
rect 62686 -112060 66158 -111348
rect 62886 -112548 66158 -112060
rect 62886 -113260 67300 -112548
rect 63086 -113748 67300 -113260
rect 63086 -114460 67500 -113748
rect 63286 -114948 67500 -114460
rect 63286 -115660 67700 -114948
rect 63600 -116148 67700 -115660
rect 63600 -116860 68842 -116148
rect 64742 -117348 68842 -116860
rect 64742 -118060 69156 -117348
rect 64942 -118548 69156 -118060
rect 64942 -119260 70298 -118548
rect 65142 -119748 70298 -119260
rect 65142 -120460 71440 -119748
rect 66284 -120948 71440 -120460
rect 66284 -121660 72582 -120948
rect 66598 -122148 72582 -121660
rect 66598 -122860 73724 -122148
rect 67740 -123348 73724 -122860
rect 67740 -124060 73924 -123348
rect -1336 -128860 2364 -124548
rect 68882 -125260 73924 -124060
rect 70024 -125748 73924 -125260
rect 70024 -126460 75066 -125748
rect 71166 -126948 75066 -126460
rect 71166 -127660 75656 -126948
rect 71366 -128148 75656 -127660
rect 71366 -129348 76430 -128148
rect 71366 -130060 77572 -129348
rect 72508 -130548 77572 -130060
rect 72508 -131260 78714 -130548
rect 73098 -131748 78714 -131260
rect 73098 -132460 79304 -131748
rect 73872 -132948 79304 -132460
rect 73872 -133660 80446 -132948
rect 75014 -134148 80446 -133660
rect 75014 -134860 80646 -134148
rect 76156 -135348 80646 -134860
rect 76156 -136060 80960 -135348
rect 76746 -136548 80960 -136060
rect 76746 -137260 82102 -136548
rect 77888 -137748 82102 -137260
rect 77888 -138460 82416 -137748
rect 78088 -138948 82416 -138460
rect 78088 -139660 82616 -138948
rect 78402 -140148 82616 -139660
rect 78402 -140860 82930 -140148
rect 79544 -141348 82930 -140860
rect 79544 -142060 84072 -141348
rect 79858 -142548 84072 -142060
rect 79858 -143260 84386 -142548
rect 80058 -143748 84386 -143260
rect 80058 -144460 84586 -143748
rect 80372 -144948 84586 -144460
rect 80372 -145660 84900 -144948
rect 81514 -146148 84900 -145660
rect 81514 -146860 85100 -146148
rect 81828 -147348 85100 -146860
rect 81828 -148060 86242 -147348
rect 82028 -148548 86242 -148060
rect 82028 -149260 87384 -148548
rect 82342 -149748 87384 -149260
rect 82342 -150460 88158 -149748
rect 82542 -150948 88158 -150460
rect 82542 -151660 88472 -150948
rect 83684 -152148 88472 -151660
rect 83684 -152860 88672 -152148
rect 84826 -153348 88672 -152860
rect 84826 -154060 89814 -153348
rect 85600 -154548 89814 -154060
rect 85600 -155260 90404 -154548
rect 85914 -155748 90404 -155260
rect 85914 -156460 91546 -155748
rect 86114 -156948 91546 -156460
rect 86114 -157660 91860 -156948
rect 87256 -158148 91860 -157660
rect 87256 -158860 93002 -158148
rect 87846 -159348 93002 -158860
rect 87846 -160060 93202 -159348
rect 88988 -160548 93202 -160060
rect 88988 -161260 93516 -160548
rect 89302 -161748 93516 -161260
rect 89302 -162460 94658 -161748
rect 90444 -162948 94658 -162460
rect 90444 -163660 95800 -162948
rect 90644 -164148 95800 -163660
rect 90644 -164860 96114 -164148
rect 90958 -166060 96114 -164860
rect 92100 -166148 96114 -166060
rect 92100 -167260 96428 -166148
rect 93242 -167348 96428 -167260
rect 93242 -168548 97202 -167348
rect 93242 -169260 98344 -168548
rect 93556 -169748 98344 -169260
rect 93556 -170460 98658 -169748
rect 93870 -170948 98658 -170460
rect 93870 -171660 99248 -170948
rect 94644 -172148 99248 -171660
rect 94644 -172860 99562 -172148
rect 95786 -173348 99562 -172860
rect 95786 -174060 100704 -173348
rect 96100 -174548 100704 -174060
rect 96100 -175260 101846 -174548
rect 96690 -175748 101846 -175260
rect 96690 -176460 102436 -175748
rect 97004 -176948 102436 -176460
rect 97004 -177660 102636 -176948
rect 98146 -178148 102636 -177660
rect 98146 -178548 102836 -178148
rect 98146 -178860 103978 -178548
rect 99288 -179748 103978 -178860
rect 99288 -180060 105120 -179748
rect 99878 -180948 105120 -180060
rect 99878 -181260 105320 -180948
rect 100078 -181348 105320 -181260
rect 100078 -181660 105520 -181348
rect 100278 -181748 105520 -181660
rect 100278 -182860 106662 -181748
rect 101420 -182948 106662 -182860
rect 101420 -184060 106862 -182948
rect 102562 -184148 106862 -184060
rect 102562 -184460 107062 -184148
rect 102762 -184860 107062 -184460
rect 102962 -185348 107062 -184860
rect 102962 -186060 107836 -185348
rect 104104 -186548 107836 -186060
rect 104104 -187260 108150 -186548
rect 104304 -188460 108150 -187260
rect 104504 -188548 108150 -188460
rect 104504 -189660 109292 -188548
rect 105278 -189748 109292 -189660
rect 105278 -190948 109492 -189748
rect 105278 -191660 110634 -190948
rect 105592 -192148 110634 -191660
rect 105592 -192860 111776 -192148
rect 106734 -193348 111776 -192860
rect 106734 -194060 111976 -193348
rect 106934 -194548 111976 -194060
rect 106934 -195260 113118 -194548
rect 108076 -195748 113118 -195260
rect 108076 -196460 114260 -195748
rect 109218 -196948 114260 -196460
rect 109218 -197660 114460 -196948
rect 109418 -198148 114460 -197660
rect 109418 -198860 115234 -198148
rect 110560 -199348 115234 -198860
rect 110560 -200060 115640 -199348
rect 111702 -200548 115640 -200060
rect 111702 -201260 116782 -200548
rect 111902 -201748 116782 -201260
rect 111902 -202460 117096 -201748
rect 112676 -202948 117096 -202460
rect 112676 -203348 117296 -202948
rect 112676 -203660 117610 -203348
rect 113082 -204548 117610 -203660
rect 113082 -204860 118752 -204548
rect 114224 -205748 118752 -204860
rect 114224 -206060 119066 -205748
rect 114538 -206460 119066 -206060
rect 114738 -206948 119066 -206460
rect 114738 -207660 120208 -206948
rect 115052 -208148 120208 -207660
rect 115052 -208860 120798 -208148
rect 116194 -209348 120798 -208860
rect 116194 -209748 120998 -209348
rect 116194 -210060 121312 -209748
rect 116508 -210948 121312 -210060
rect 116508 -211260 121626 -210948
rect 117650 -212148 121626 -211260
rect 117650 -212460 121826 -212148
rect 118240 -212548 121826 -212460
rect 118240 -212860 122140 -212548
rect 118440 -213748 122140 -212860
rect 118440 -214060 122730 -213748
rect 118754 -214948 122730 -214060
rect 118754 -215260 123044 -214948
rect 119068 -215660 123044 -215260
rect 119268 -216148 123044 -215660
rect 119268 -216860 123634 -216148
rect 119582 -217348 123634 -216860
rect 119582 -218060 123948 -217348
rect 120172 -218548 123948 -218060
rect 120172 -219260 125090 -218548
rect 120486 -219748 125090 -219260
rect 120486 -220148 125290 -219748
rect 120486 -220460 125604 -220148
rect 121076 -221348 125604 -220460
rect 121076 -221660 125918 -221348
rect 121390 -222548 125918 -221660
rect 121390 -222860 126232 -222548
rect 122532 -223260 126232 -222860
rect 122732 -223748 126232 -223260
rect 122732 -224460 126546 -223748
rect 123046 -224948 126546 -224460
rect 123046 -225660 127688 -224948
rect 123360 -226148 127688 -225660
rect 123360 -226860 128278 -226148
rect 123674 -228060 128278 -226860
rect 123988 -228148 128278 -228060
rect 123988 -229260 129420 -228148
rect 125130 -229348 129420 -229260
rect 125130 -230548 129734 -229348
rect 125130 -231260 129934 -230548
rect 125720 -231748 129934 -231260
rect 125720 -232460 130248 -231748
rect 126862 -232948 130248 -232460
rect 126862 -233660 130448 -232948
rect 127176 -234148 130448 -233660
rect 127176 -234860 130648 -234148
rect 127376 -235348 130648 -234860
rect 127376 -236060 130848 -235348
rect 127690 -236548 130848 -236060
rect 127690 -237260 131162 -236548
rect 127890 -237748 131162 -237260
rect 127890 -238460 132304 -237748
rect 128090 -238948 132304 -238460
rect 128090 -239660 132504 -238948
rect 128290 -240148 132504 -239660
rect 128290 -240860 132704 -240148
rect 128604 -241348 132704 -240860
rect 128604 -242060 133846 -241348
rect 129746 -242548 133846 -242060
rect 129746 -243260 134160 -242548
rect 129946 -243748 134160 -243260
rect 129946 -244460 135302 -243748
rect 130146 -244948 135302 -244460
rect 130146 -245660 136444 -244948
rect 131288 -246148 136444 -245660
rect 131288 -246860 137586 -246148
rect 131602 -247348 137586 -246860
rect 131602 -248060 138728 -247348
rect 132744 -248548 138728 -248060
rect 132744 -249260 138928 -248548
rect 133886 -250460 138928 -249260
rect 135028 -251660 138928 -250460
rect 136170 -252860 138928 -251660
<< viali >>
rect 5457 8925 5491 8959
rect 5273 8789 5307 8823
rect 4445 3009 4479 3043
rect 4353 2805 4387 2839
rect 1777 2397 1811 2431
rect 1409 2329 1443 2363
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8956 5503 8959
rect 6454 8956 6460 8968
rect 5491 8928 6460 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 5258 3136 5264 3188
rect 5316 3136 5322 3188
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 5276 3040 5304 3136
rect 4479 3012 5304 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4338 2796 4344 2848
rect 4396 2796 4402 2848
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 4338 2428 4344 2440
rect 1811 2400 4344 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6460 8916 6512 8968
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 5264 3136 5316 3188
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 4344 2388 4396 2440
rect 20 2320 72 2372
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 6458 10624 6514 11424
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 6472 8974 6500 10624
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 5276 3194 5304 8774
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 4356 2446 4384 2790
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 18 0 74 800
<< via2 >>
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
<< metal3 >>
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__inv_2  _0_
timestamp 1758435568
transform -1 0 4508 0 -1 3264
box -38 -2000 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 1758435568
transform 1 0 1932 0 1 2176
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 1758435568
transform 1 0 3036 0 1 2176
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1758435568
transform 1 0 3588 0 1 2176
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1758435568
transform 1 0 3772 0 1 2176
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_41
timestamp 1758435568
transform 1 0 4876 0 1 2176
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_47
timestamp 1758435568
transform 1 0 5428 0 1 2176
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1758435568
transform 1 0 1380 0 -1 3264
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1758435568
transform 1 0 2484 0 -1 3264
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27
timestamp 1758435568
transform 1 0 3588 0 -1 3264
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_33
timestamp 1758435568
transform 1 0 4140 0 -1 3264
box -38 -1200 200 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_37
timestamp 1758435568
transform 1 0 4508 0 -1 3264
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_45
timestamp 1758435568
transform 1 0 5244 0 -1 3264
box -38 -1200 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1758435568
transform 1 0 1380 0 1 3264
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1758435568
transform 1 0 2484 0 1 3264
box -38 -1200 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1758435568
transform 1 0 3588 0 1 3264
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1758435568
transform 1 0 3772 0 1 3264
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 1758435568
transform 1 0 4876 0 1 3264
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 1758435568
transform 1 0 5428 0 1 3264
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1758435568
transform 1 0 1380 0 -1 4352
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1758435568
transform 1 0 2484 0 -1 4352
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1758435568
transform 1 0 3588 0 -1 4352
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_39
timestamp 1758435568
transform 1 0 4692 0 -1 4352
box -38 -1200 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_47
timestamp 1758435568
transform 1 0 5428 0 -1 4352
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1758435568
transform 1 0 1380 0 1 4352
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1758435568
transform 1 0 2484 0 1 4352
box -38 -1200 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1758435568
transform 1 0 3588 0 1 4352
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1758435568
transform 1 0 3772 0 1 4352
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 1758435568
transform 1 0 4876 0 1 4352
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 1758435568
transform 1 0 5428 0 1 4352
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1758435568
transform 1 0 1380 0 -1 5440
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1758435568
transform 1 0 2484 0 -1 5440
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1758435568
transform 1 0 3588 0 -1 5440
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_39
timestamp 1758435568
transform 1 0 4692 0 -1 5440
box -38 -1200 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_47
timestamp 1758435568
transform 1 0 5428 0 -1 5440
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1758435568
transform 1 0 1380 0 1 5440
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1758435568
transform 1 0 2484 0 1 5440
box -38 -1200 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1758435568
transform 1 0 3588 0 1 5440
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1758435568
transform 1 0 3772 0 1 5440
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 1758435568
transform 1 0 4876 0 1 5440
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 1758435568
transform 1 0 5428 0 1 5440
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1758435568
transform 1 0 1380 0 -1 6528
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1758435568
transform 1 0 2484 0 -1 6528
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1758435568
transform 1 0 3588 0 -1 6528
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 1758435568
transform 1 0 4692 0 -1 6528
box -38 -1200 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_47
timestamp 1758435568
transform 1 0 5428 0 -1 6528
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1758435568
transform 1 0 1380 0 1 6528
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1758435568
transform 1 0 2484 0 1 6528
box -38 -1200 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1758435568
transform 1 0 3588 0 1 6528
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1758435568
transform 1 0 3772 0 1 6528
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 1758435568
transform 1 0 4876 0 1 6528
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_47
timestamp 1758435568
transform 1 0 5428 0 1 6528
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1758435568
transform 1 0 1380 0 -1 7616
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1758435568
transform 1 0 2484 0 -1 7616
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1758435568
transform 1 0 3588 0 -1 7616
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 1758435568
transform 1 0 4692 0 -1 7616
box -38 -1200 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 1758435568
transform 1 0 5428 0 -1 7616
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1758435568
transform 1 0 1380 0 1 7616
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1758435568
transform 1 0 2484 0 1 7616
box -38 -1200 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1758435568
transform 1 0 3588 0 1 7616
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1758435568
transform 1 0 3772 0 1 7616
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_41
timestamp 1758435568
transform 1 0 4876 0 1 7616
box -38 -1200 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_47
timestamp 1758435568
transform 1 0 5428 0 1 7616
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1758435568
transform 1 0 1380 0 -1 8704
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1758435568
transform 1 0 2484 0 -1 8704
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1758435568
transform 1 0 3588 0 -1 8704
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_39
timestamp 1758435568
transform 1 0 4692 0 -1 8704
box -38 -1200 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_47
timestamp 1758435568
transform 1 0 5428 0 -1 8704
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1758435568
transform 1 0 1380 0 1 8704
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1758435568
transform 1 0 2484 0 1 8704
box -38 -1200 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1758435568
transform 1 0 3588 0 1 8704
box -38 -1200 200 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1758435568
transform 1 0 3772 0 1 8704
box -38 -1200 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_41
timestamp 1758435568
transform 1 0 4876 0 1 8704
box -38 -1200 406 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1758435568
transform -1 0 5520 0 1 8704
box -38 -2000 314 592
use sky130_fd_sc_hd__clkbuf_4  output2
timestamp 1758435568
transform -1 0 1932 0 1 2176
box -38 -2000 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1758435568
transform 1 0 1104 0 1 2176
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1758435568
transform -1 0 5796 0 1 2176
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1758435568
transform 1 0 1104 0 -1 3264
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1758435568
transform -1 0 5796 0 -1 3264
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1758435568
transform 1 0 1104 0 1 3264
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1758435568
transform -1 0 5796 0 1 3264
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1758435568
transform 1 0 1104 0 -1 4352
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1758435568
transform -1 0 5796 0 -1 4352
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1758435568
transform 1 0 1104 0 1 4352
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1758435568
transform -1 0 5796 0 1 4352
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1758435568
transform 1 0 1104 0 -1 5440
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1758435568
transform -1 0 5796 0 -1 5440
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1758435568
transform 1 0 1104 0 1 5440
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1758435568
transform -1 0 5796 0 1 5440
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1758435568
transform 1 0 1104 0 -1 6528
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1758435568
transform -1 0 5796 0 -1 6528
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1758435568
transform 1 0 1104 0 1 6528
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1758435568
transform -1 0 5796 0 1 6528
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1758435568
transform 1 0 1104 0 -1 7616
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1758435568
transform -1 0 5796 0 -1 7616
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1758435568
transform 1 0 1104 0 1 7616
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1758435568
transform -1 0 5796 0 1 7616
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1758435568
transform 1 0 1104 0 -1 8704
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1758435568
transform -1 0 5796 0 -1 8704
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1758435568
transform 1 0 1104 0 1 8704
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1758435568
transform -1 0 5796 0 1 8704
box -38 -1200 314 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_0
timestamp 1758435568
transform 1 0 6518 0 1 -1200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_1
timestamp 1758435568
transform 1 0 7660 0 1 -2400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_2
timestamp 1758435568
transform 1 0 10166 0 1 -6000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_3
timestamp 1758435568
transform 1 0 11308 0 1 -7200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_4
timestamp 1758435568
transform 1 0 13040 0 1 -9600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_5
timestamp 1758435568
transform 1 0 14696 0 1 -13200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_6
timestamp 1758435568
transform 1 0 16666 0 1 -18000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_7
timestamp 1758435568
transform 1 0 18836 0 1 -24000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_8
timestamp 1758435568
transform 1 0 19978 0 1 -25200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_9
timestamp 1758435568
transform 1 0 22408 0 1 -30000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_10
timestamp 1758435568
transform 1 0 24140 0 1 -32400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_11
timestamp 1758435568
transform 1 0 25596 0 1 -34800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_12
timestamp 1758435568
transform 1 0 27252 0 1 -38400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_13
timestamp 1758435568
transform 1 0 28394 0 1 -39600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_14
timestamp 1758435568
transform 1 0 30938 0 1 -45200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_15
timestamp 1758435568
transform 1 0 33298 0 1 -50000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_16
timestamp 1758435568
transform 1 0 34440 0 1 -51200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_17
timestamp 1758435568
transform 1 0 36572 0 1 -55200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_18
timestamp 1758435568
transform 1 0 37714 0 1 -56400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_19
timestamp 1758435568
transform 1 0 39256 0 1 -58400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_20
timestamp 1758435568
transform 1 0 41886 0 1 -65200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_21
timestamp 1758435568
transform 1 0 43228 0 1 -67600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_22
timestamp 1758435568
transform 1 0 44370 0 1 -68800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_23
timestamp 1758435568
transform 1 0 45712 0 1 -71200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_24
timestamp 1758435568
transform 1 0 46854 0 1 -72400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_25
timestamp 1758435568
transform 1 0 49376 0 1 -77200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_26
timestamp 1758435568
transform 1 0 51346 0 1 -81200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_27
timestamp 1758435568
transform 1 0 52802 0 1 -83600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_28
timestamp 1758435568
transform 1 0 57684 0 1 -95200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_29
timestamp 1758435568
transform 1 0 60282 0 1 -101600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_30
timestamp 1758435568
transform 1 0 62014 0 1 -104800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_31
timestamp 1758435568
transform 1 0 64898 0 1 -114400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_32
timestamp 1758435568
transform 1 0 66440 0 1 -118000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_33
timestamp 1758435568
transform 1 0 67896 0 1 -120400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_34
timestamp 1758435568
transform 1 0 69038 0 1 -121600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_35
timestamp 1758435568
transform 1 0 70180 0 1 -122800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_36
timestamp 1758435568
transform 1 0 71322 0 1 -124000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_37
timestamp 1758435568
transform 1 0 -38 0 1 -126400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_38
timestamp 1758435568
transform 1 0 72664 0 1 -127600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_39
timestamp 1758435568
transform 1 0 75170 0 1 -131200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_40
timestamp 1758435568
transform 1 0 76312 0 1 -132400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_41
timestamp 1758435568
transform 1 0 78044 0 1 -134800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_42
timestamp 1758435568
transform 1 0 79700 0 1 -138400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_43
timestamp 1758435568
transform 1 0 81670 0 1 -143200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_44
timestamp 1758435568
transform 1 0 83840 0 1 -149200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_45
timestamp 1758435568
transform 1 0 84982 0 1 -150400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_46
timestamp 1758435568
transform 1 0 87412 0 1 -155200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_47
timestamp 1758435568
transform 1 0 89144 0 1 -157600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_48
timestamp 1758435568
transform 1 0 90600 0 1 -160000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_49
timestamp 1758435568
transform 1 0 92256 0 1 -163600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_50
timestamp 1758435568
transform 1 0 93398 0 1 -164800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_51
timestamp 1758435568
transform 1 0 95942 0 1 -170400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_52
timestamp 1758435568
transform 1 0 98302 0 1 -175200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_53
timestamp 1758435568
transform 1 0 99444 0 1 -176400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_54
timestamp 1758435568
transform 1 0 101576 0 1 -180400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_55
timestamp 1758435568
transform 1 0 102718 0 1 -181600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_56
timestamp 1758435568
transform 1 0 104260 0 1 -183600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_57
timestamp 1758435568
transform 1 0 106890 0 1 -190400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_58
timestamp 1758435568
transform 1 0 108232 0 1 -192800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_59
timestamp 1758435568
transform 1 0 109374 0 1 -194000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_60
timestamp 1758435568
transform 1 0 110716 0 1 -196400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_61
timestamp 1758435568
transform 1 0 111858 0 1 -197600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_62
timestamp 1758435568
transform 1 0 114380 0 1 -202400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_63
timestamp 1758435568
transform 1 0 116350 0 1 -206400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_64
timestamp 1758435568
transform 1 0 117806 0 1 -208800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_65
timestamp 1758435568
transform 1 0 122688 0 1 -220400
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_66
timestamp 1758435568
transform 1 0 125286 0 1 -226800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_67
timestamp 1758435568
transform 1 0 127018 0 1 -230000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_68
timestamp 1758435568
transform 1 0 129902 0 1 -239600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_69
timestamp 1758435568
transform 1 0 131444 0 1 -243200
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_70
timestamp 1758435568
transform 1 0 132900 0 1 -245600
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_71
timestamp 1758435568
transform 1 0 134042 0 1 -246800
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_72
timestamp 1758435568
transform 1 0 135184 0 1 -248000
box -38 -1200 1142 592
use sky130_ef_sc_hd__decap_12  sky130_ef_sc_hd__decap_12_73
timestamp 1758435568
transform 1 0 136326 0 1 -249200
box -38 -1200 1142 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0
timestamp 1758435568
transform 1 0 29536 0 1 -40800
box -38 -2000 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_1
timestamp 1758435568
transform 1 0 94540 0 1 -166000
box -38 -2000 314 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_0
timestamp 1758435568
transform 1 0 61424 0 1 -102800
box -38 -2000 590 592
use sky130_fd_sc_hd__clkbuf_4  sky130_fd_sc_hd__clkbuf_4_1
timestamp 1758435568
transform 1 0 126428 0 1 -228000
box -38 -2000 590 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_0
timestamp 1758435568
transform 1 0 14382 0 1 -12000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_1
timestamp 1758435568
transform 1 0 15838 0 1 -14400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_2
timestamp 1758435568
transform 1 0 16352 0 1 -16800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_3
timestamp 1758435568
transform 1 0 17808 0 1 -19200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_4
timestamp 1758435568
transform 1 0 18322 0 1 -21600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_5
timestamp 1758435568
transform 1 0 21894 0 1 -27600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_6
timestamp 1758435568
transform 1 0 25282 0 1 -33600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_7
timestamp 1758435568
transform 1 0 26938 0 1 -37200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_8
timestamp 1758435568
transform 1 0 29850 0 1 -42800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_9
timestamp 1758435568
transform 1 0 32080 0 1 -46400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_10
timestamp 1758435568
transform 1 0 32984 0 1 -48800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_11
timestamp 1758435568
transform 1 0 50518 0 1 -78400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_12
timestamp 1758435568
transform 1 0 51032 0 1 -80000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_13
timestamp 1758435568
transform 1 0 52488 0 1 -82400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_14
timestamp 1758435568
transform 1 0 54734 0 1 -86400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_15
timestamp 1758435568
transform 1 0 55048 0 1 -87600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_16
timestamp 1758435568
transform 1 0 55562 0 1 -89200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_17
timestamp 1758435568
transform 1 0 56466 0 1 -91600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_18
timestamp 1758435568
transform 1 0 57370 0 1 -94000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_19
timestamp 1758435568
transform 1 0 59026 0 1 -96800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_20
timestamp 1758435568
transform 1 0 59340 0 1 -98000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_21
timestamp 1758435568
transform 1 0 59654 0 1 -99200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_22
timestamp 1758435568
transform 1 0 59968 0 1 -100400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_23
timestamp 1758435568
transform 1 0 63156 0 1 -106000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_24
timestamp 1758435568
transform 1 0 63670 0 1 -108400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_25
timestamp 1758435568
transform 1 0 64584 0 1 -113200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_26
timestamp 1758435568
transform 1 0 67582 0 1 -119200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_27
timestamp 1758435568
transform 1 0 79386 0 1 -137200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_28
timestamp 1758435568
transform 1 0 80842 0 1 -139600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_29
timestamp 1758435568
transform 1 0 81356 0 1 -142000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_30
timestamp 1758435568
transform 1 0 82812 0 1 -144400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_31
timestamp 1758435568
transform 1 0 83326 0 1 -146800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_32
timestamp 1758435568
transform 1 0 86898 0 1 -152800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_33
timestamp 1758435568
transform 1 0 90286 0 1 -158800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_34
timestamp 1758435568
transform 1 0 91942 0 1 -162400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_35
timestamp 1758435568
transform 1 0 94854 0 1 -168000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_36
timestamp 1758435568
transform 1 0 97084 0 1 -171600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_37
timestamp 1758435568
transform 1 0 97988 0 1 -174000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_38
timestamp 1758435568
transform 1 0 115522 0 1 -203600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_39
timestamp 1758435568
transform 1 0 116036 0 1 -205200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_40
timestamp 1758435568
transform 1 0 117492 0 1 -207600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_41
timestamp 1758435568
transform 1 0 119738 0 1 -211600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_42
timestamp 1758435568
transform 1 0 120052 0 1 -212800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_43
timestamp 1758435568
transform 1 0 120566 0 1 -214400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_44
timestamp 1758435568
transform 1 0 121470 0 1 -216800
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_45
timestamp 1758435568
transform 1 0 122374 0 1 -219200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_46
timestamp 1758435568
transform 1 0 124030 0 1 -222000
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_47
timestamp 1758435568
transform 1 0 124344 0 1 -223200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_48
timestamp 1758435568
transform 1 0 124658 0 1 -224400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_49
timestamp 1758435568
transform 1 0 124972 0 1 -225600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_50
timestamp 1758435568
transform 1 0 128160 0 1 -231200
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_51
timestamp 1758435568
transform 1 0 128674 0 1 -233600
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_52
timestamp 1758435568
transform 1 0 129588 0 1 -238400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_3  sky130_fd_sc_hd__decap_3_53
timestamp 1758435568
transform 1 0 132586 0 1 -244400
box -38 -1200 314 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_0
timestamp 1758435568
transform 1 0 48970 0 1 -76000
box -38 -1200 406 592
use sky130_fd_sc_hd__decap_4  sky130_fd_sc_hd__decap_4_1
timestamp 1758435568
transform 1 0 113974 0 1 -201200
box -38 -1200 406 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_0
timestamp 1758435568
transform 1 0 8802 0 1 -3600
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_1
timestamp 1758435568
transform 1 0 12450 0 1 -8400
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_2
timestamp 1758435568
transform 1 0 23550 0 1 -31200
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_3
timestamp 1758435568
transform 1 0 32394 0 1 -47600
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_4
timestamp 1758435568
transform 1 0 35582 0 1 -52400
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_5
timestamp 1758435568
transform 1 0 53944 0 1 -84800
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_6
timestamp 1758435568
transform 1 0 55876 0 1 -90400
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_7
timestamp 1758435568
transform 1 0 56780 0 1 -92800
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_8
timestamp 1758435568
transform 1 0 73806 0 1 -128800
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_9
timestamp 1758435568
transform 1 0 77454 0 1 -133600
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_10
timestamp 1758435568
transform 1 0 88554 0 1 -156400
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_11
timestamp 1758435568
transform 1 0 97398 0 1 -172800
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_12
timestamp 1758435568
transform 1 0 100586 0 1 -177600
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_13
timestamp 1758435568
transform 1 0 118948 0 1 -210000
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_14
timestamp 1758435568
transform 1 0 120880 0 1 -215600
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_6  sky130_fd_sc_hd__decap_6_15
timestamp 1758435568
transform 1 0 121784 0 1 -218000
box -38 -1200 590 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_0
timestamp 1758435568
transform 1 0 0 0 1 600
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_1
timestamp 1758435568
transform 1 0 9392 0 1 -4800
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_2
timestamp 1758435568
transform 1 0 21120 0 1 -26400
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_3
timestamp 1758435568
transform 1 0 30164 0 1 -44000
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_4
timestamp 1758435568
transform 1 0 40798 0 1 -62000
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_5
timestamp 1758435568
transform 1 0 48196 0 1 -74800
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_6
timestamp 1758435568
transform 1 0 74396 0 1 -130000
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_7
timestamp 1758435568
transform 1 0 86124 0 1 -151600
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_8
timestamp 1758435568
transform 1 0 95168 0 1 -169200
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_9
timestamp 1758435568
transform 1 0 105802 0 1 -187200
box -38 -1200 774 592
use sky130_fd_sc_hd__decap_8  sky130_fd_sc_hd__decap_8_10
timestamp 1758435568
transform 1 0 113200 0 1 -200000
box -38 -1200 774 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0
timestamp 1758435568
transform 1 0 14182 0 1 -10800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1758435568
transform 1 0 16152 0 1 -15600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1758435568
transform 1 0 18122 0 1 -20400
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1758435568
transform 1 0 18636 0 1 -22800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1758435568
transform 1 0 22208 0 1 -28800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1758435568
transform 1 0 26738 0 1 -36000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1758435568
transform 1 0 36172 0 1 -53600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1758435568
transform 1 0 40398 0 1 -59600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1758435568
transform 1 0 40598 0 1 -60800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1758435568
transform 1 0 43028 0 1 -66400
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1758435568
transform 1 0 45512 0 1 -70000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1758435568
transform 1 0 47996 0 1 -73600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1758435568
transform 1 0 63470 0 1 -107200
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1758435568
transform 1 0 63984 0 1 -109600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1758435568
transform 1 0 64184 0 1 -110800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1758435568
transform 1 0 64384 0 1 -112000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1758435568
transform 1 0 66040 0 1 -115600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1758435568
transform 1 0 66240 0 1 -116800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1758435568
transform 1 0 72464 0 1 -125200
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1758435568
transform 1 0 79186 0 1 -136000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1758435568
transform 1 0 81156 0 1 -140800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21
timestamp 1758435568
transform 1 0 83126 0 1 -145600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_22
timestamp 1758435568
transform 1 0 83640 0 1 -148000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_23
timestamp 1758435568
transform 1 0 87212 0 1 -154000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_24
timestamp 1758435568
transform 1 0 91742 0 1 -161200
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_25
timestamp 1758435568
transform 1 0 101176 0 1 -178800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_26
timestamp 1758435568
transform 1 0 105402 0 1 -184800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_27
timestamp 1758435568
transform 1 0 105602 0 1 -186000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_28
timestamp 1758435568
transform 1 0 108032 0 1 -191600
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_29
timestamp 1758435568
transform 1 0 110516 0 1 -195200
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_30
timestamp 1758435568
transform 1 0 113000 0 1 -198800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_31
timestamp 1758435568
transform 1 0 128474 0 1 -232400
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_32
timestamp 1758435568
transform 1 0 128988 0 1 -234800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_33
timestamp 1758435568
transform 1 0 129188 0 1 -236000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_34
timestamp 1758435568
transform 1 0 129388 0 1 -237200
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_35
timestamp 1758435568
transform 1 0 131044 0 1 -240800
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_36
timestamp 1758435568
transform 1 0 131244 0 1 -242000
box -38 -1200 200 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_37
timestamp 1758435568
transform 1 0 137468 0 1 -250400
box -38 -1200 200 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_0
timestamp 1758435568
transform 1 0 41572 0 1 -63200
box -38 -2000 314 592
use sky130_fd_sc_hd__inv_2  sky130_fd_sc_hd__inv_2_1
timestamp 1758435568
transform 1 0 106576 0 1 -188400
box -38 -2000 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1758435568
transform 1 0 36372 0 1 -54800
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1758435568
transform 1 0 38856 0 1 -57600
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1758435568
transform 1 0 39056 0 1 -58000
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1758435568
transform 1 0 50832 0 1 -79600
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1758435568
transform 1 0 54534 0 1 -86000
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1758435568
transform 1 0 55362 0 1 -88800
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1758435568
transform 1 0 58826 0 1 -96400
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1758435568
transform 1 0 101376 0 1 -180000
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_8
timestamp 1758435568
transform 1 0 103860 0 1 -182800
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_9
timestamp 1758435568
transform 1 0 104060 0 1 -183200
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_10
timestamp 1758435568
transform 1 0 115836 0 1 -204800
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_11
timestamp 1758435568
transform 1 0 119538 0 1 -211200
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_12
timestamp 1758435568
transform 1 0 120366 0 1 -214000
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_13
timestamp 1758435568
transform 1 0 123830 0 1 -221600
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1758435568
transform 1 0 3680 0 1 2176
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1758435568
transform 1 0 3680 0 1 3264
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1758435568
transform 1 0 3680 0 1 4352
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1758435568
transform 1 0 3680 0 1 5440
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1758435568
transform 1 0 3680 0 1 6528
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1758435568
transform 1 0 3680 0 1 7616
box -38 -400 200 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1758435568
transform 1 0 3680 0 1 8704
box -38 -400 200 592
<< labels >>
rlabel metal1 s 3450 8704 3450 8704 4 VGND
rlabel metal1 s 3450 9248 3450 9248 4 VPWR
rlabel metal1 s 5980 8942 5980 8942 4 in
rlabel metal1 s 4876 3026 4876 3026 4 net1
rlabel metal1 s 3082 2414 3082 2414 4 net2
rlabel metal2 s 46 1554 46 1554 4 out
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 6458 10624 6514 11424 0 FreeSans 280 90 0 0 in
port 3 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 out
port 4 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VGND
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VPWR
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 in
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 out
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
