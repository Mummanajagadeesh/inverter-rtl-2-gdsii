magic
tech sky130A
magscale 1 2
timestamp 1758368339
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37584
<< metal2 >>
rect 39302 39200 39358 40000
rect 18 0 74 800
<< obsm2 >>
rect 20 39144 39246 39200
rect 20 856 39356 39144
rect 130 800 39356 856
<< obsm3 >>
rect 4210 2143 35906 37569
<< metal4 >>
rect 4208 2128 4528 37584
rect 4868 2128 5188 37584
rect 34928 2128 35248 37584
rect 35588 2128 35908 37584
<< metal5 >>
rect 1056 36642 38872 36962
rect 1056 35982 38872 36302
rect 1056 6006 38872 6326
rect 1056 5346 38872 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 38872 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 38872 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 38872 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 38872 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 39302 39200 39358 40000 6 in
port 3 nsew signal input
rlabel metal2 s 18 0 74 800 6 out
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 445846
string GDS_FILE /openlane/designs/inverter/runs/myrun/results/signoff/inverter.magic.gds
string GDS_START 34008
<< end >>

