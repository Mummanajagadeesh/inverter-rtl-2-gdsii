magic
tech sky130A
magscale 1 2
timestamp 1758433797
<< checkpaint >>
rect -3918 -3932 10450 15356
<< viali >>
rect 5457 8925 5491 8959
rect 5273 8789 5307 8823
rect 4445 3009 4479 3043
rect 4353 2805 4387 2839
rect 1777 2397 1811 2431
rect 1409 2329 1443 2363
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8956 5503 8959
rect 6454 8956 6460 8968
rect 5491 8928 6460 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 5258 3136 5264 3188
rect 5316 3136 5322 3188
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 5276 3040 5304 3136
rect 4479 3012 5304 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4338 2796 4344 2848
rect 4396 2796 4402 2848
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1765 2431 1823 2437
rect 1765 2397 1777 2431
rect 1811 2428 1823 2431
rect 4338 2428 4344 2440
rect 1811 2400 4344 2428
rect 1811 2397 1823 2400
rect 1765 2391 1823 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 6460 8916 6512 8968
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 5264 3136 5316 3188
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 4344 2388 4396 2440
rect 20 2320 72 2372
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 6458 10624 6514 11424
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 6472 8974 6500 10624
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 5276 3194 5304 8774
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 4356 2446 4384 2790
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 32 800 60 2314
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 18 0 74 800
<< via2 >>
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
<< metal3 >>
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__inv_2  _0_
timestamp 0
transform -1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9
timestamp 0
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21
timestamp 0
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_47
timestamp 0
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_33
timestamp 0
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_37
timestamp 0
transform 1 0 4508 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_45
timestamp 0
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_47
timestamp 0
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_47
timestamp 0
transform 1 0 5428 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 0
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_47
timestamp 0
transform 1 0 5428 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_47
timestamp 0
transform 1 0 5428 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_47
timestamp 0
transform 1 0 5428 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_47
timestamp 0
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 0
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_47
timestamp 0
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_47
timestamp 0
transform 1 0 5428 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform -1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output2
timestamp 0
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
rlabel metal1 s 3450 8704 3450 8704 4 VGND
rlabel metal1 s 3450 9248 3450 9248 4 VPWR
rlabel metal1 s 5980 8942 5980 8942 4 in
rlabel metal1 s 4876 3026 4876 3026 4 net1
rlabel metal1 s 3082 2414 3082 2414 4 net2
rlabel metal2 s 46 1554 46 1554 4 out
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal2 s 6458 10624 6514 11424 0 FreeSans 280 90 0 0 in
port 3 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 out
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
